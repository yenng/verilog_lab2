module download(
	input [9:0] SW,								//IR and Enter is the control signal.
	input [0:0] KEY,							//Aeq0 and Apos is value of part of PCload.
	output [9:0] LEDR,													//status signal
	output [3:0] LEDG											//state
	);
	
	controlUnit	try(SW[9:7],SW[6],SW[5],SW[4],KEY[0],SW[0],LEDR[9],LEDR[8],LEDR[7],LEDR[6],LEDR[5],LEDR[4],LEDR[3],LEDR[2],LEDR[1:0],LEDG[3:0]);
	
endmodule