module controlUnit(
	input [2:0] IR,								//IR and Enter is the control signal.
	input Enter, Aeq0, Apos, clock, reset,		//Aeq0 and Apos is value of part of PCload.
	output reg IRload, JMPmux, PCload, Meminst, MemWr, Aload, Sub, Halt,	//status signal
	output reg [1:0] Asel,													//status signal
	output reg [3:0] state													//state
	);
	
	reg [3:0] nextstate;
	parameter start = 0, fetch = 1, decode = 2, load = 8, store = 9, add = 10, sub = 11, Input = 12, jz = 13, jpos = 14, halt = 15;
	
	always@(posedge clock, posedge reset) 	//Control the changing of state by using clock.
	begin
		if(reset)
			state <= start;					//If reset = 1, the state changes to start.
		else
			state <= nextstate;
	end
	
	always@(IR,Enter,state,Apos,Aeq0)  
	begin      
		case(state)
			start:	begin
				{IRload, JMPmux, PCload, Meminst, MemWr, Asel, Aload, Sub, Halt} = 10'b 0000000000;
				nextstate = fetch;
				end
			fetch:	begin
				{IRload, JMPmux, PCload, Meminst, MemWr, Asel, Aload, Sub, Halt} = 10'b 1010000000;
				nextstate = decode;
				end
			decode:	begin
				{IRload, JMPmux, PCload, Meminst, MemWr, Asel, Aload, Sub, Halt} = 10'b 0001000000;
				case(IR)								//NextState of this state depend on control signal IR.
					3'b 000: nextstate = load;
					3'b 001: nextstate = store;
					3'b 010: nextstate = add;
					3'b 011: nextstate = sub;
					3'b 100: nextstate = Input;
					3'b 101: nextstate = jz;
					3'b 110: nextstate = jpos;
					3'b 111: nextstate = halt;
					default: nextstate = decode;
				endcase
				end
			load:	begin
				{IRload, JMPmux, PCload, Meminst, MemWr, Asel, Aload, Sub, Halt} = 10'b 0000010100; 
				nextstate = start;
				end
			store:	begin
				{IRload, JMPmux, PCload, Meminst, MemWr, Asel, Aload, Sub, Halt} = 10'b 0001100000;
				nextstate = start;
				end
			add:	begin
				{IRload, JMPmux, PCload, Meminst, MemWr, Asel, Aload, Sub, Halt} = 10'b 0000000100;
				nextstate = start;
				end
			sub:	begin
				{IRload, JMPmux, PCload, Meminst, MemWr, Asel, Aload, Sub, Halt} = 10'b 0000000110;
				nextstate = start;
				end
			Input:	begin
				{IRload, JMPmux, PCload, Meminst, MemWr, Asel, Aload, Sub, Halt} = 10'b 0000001100;
				if(Enter)							//NextState of this state depend on control signal Enter.
					nextstate = start;
				else
					nextstate = Input;
				end
			jz:		begin
				{IRload, JMPmux, Meminst, MemWr, Asel, Aload, Sub, Halt} = 9'b 010000000;
				PCload = Aeq0;						//If A equal to zero, PCload = 1.
				nextstate = start;	
				end
			jpos:	begin
				{IRload, JMPmux, Meminst, MemWr, Asel, Aload, Sub, Halt} = 9'b 010000000;
				PCload = Apos;						//If A is positive, PCload = 1.
				nextstate = start;
				end
			halt:	begin
				{IRload, JMPmux, PCload, Meminst, MemWr, Asel, Aload, Sub, Halt} = 10'b 0000000001;
				nextstate = halt;
				end
			default:begin
				{IRload, JMPmux, PCload, Meminst, MemWr, Asel, Aload, Sub, Halt} = 10'b 0000000000;
				nextstate = fetch;
				end
		endcase
	end
//	assign displayState = state;
endmodule 